LIBRARY IEEE;
LIBRARY WORK;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
ENTITY SRAM IS
  PORT (
    CLOCK : IN STD_LOGIC;
    IO_WRITE : IN STD_LOGIC;
    SRAM_UPPER_ADDR : IN STD_LOGIC;
    SRAM_LOWER_ADDR : IN STD_LOGIC;
    SRAM_DATA : IN STD_LOGIC;
    SRAM_INC_DATA : IN STD_LOGIC;
    SRAM_ADDR_JPOS : IN STD_LOGIC;
    SRAM_ADDR_JNEG : IN STD_LOGIC;
    IO_DATA : INOUT STD_LOGIC_VECTOR(15 DOWNTO 0);
    SRAM_CE_N : OUT STD_LOGIC;
    SRAM_WE_N : OUT STD_LOGIC;
    SRAM_OE_N : OUT STD_LOGIC;
    SRAM_UB_N : OUT STD_LOGIC;
    SRAM_LB_N : OUT STD_LOGIC;
    SRAM_ADDR : OUT STD_LOGIC_VECTOR(17 DOWNTO 0)
  );
END SRAM;

ARCHITECTURE bdf_type OF SRAM IS
  TYPE STATE_TYPE IS (
    IDLE,
    READ_UPPER,
    WRITE_UPPER,
    READ_LOWER,
    WRITE_LOWER,
    SRAM_READ,
    SRAM_INC_READ,
    SRAM_WRITE,
    SRAM_INC_WRITE,
    JUMP_POS,
    JUMP_NEG
  );
  SIGNAL PREV_STATE : STATE_TYPE;
  SIGNAL STATE : STATE_TYPE;
  SIGNAL SRAM_ADDR_ALTERA_SYNTHESIZED : STD_LOGIC_VECTOR(17 DOWNTO 0) := "000000000000000000";

BEGIN
  SRAM_ADDR <= SRAM_ADDR_ALTERA_SYNTHESIZED;
  SRAM_CE_N <= '0';
  SRAM_UB_N <= '0';
  SRAM_LB_N <= '0';
  
  PROCESS (CLOCK)
  BEGIN
    IF (RISING_EDGE(CLOCK)) THEN
    
		IF (SRAM_UPPER_ADDR = '1' AND IO_WRITE = '0') THEN
			STATE <= READ_UPPER;
		ELSIF (SRAM_UPPER_ADDR = '1' AND IO_WRITE = '1') THEN
			STATE <= WRITE_UPPER;
		ELSIF (SRAM_LOWER_ADDR = '1' AND IO_WRITE = '0') THEN
			STATE <= READ_LOWER;
		ELSIF (SRAM_LOWER_ADDR = '1' AND IO_WRITE = '1') THEN
			STATE <= WRITE_LOWER;
		ELSIF (SRAM_DATA = '1' AND IO_WRITE = '0') THEN
			STATE <= SRAM_READ;
		ELSIF (SRAM_INC_DATA = '1' AND IO_WRITE = '0') THEN
			STATE <= SRAM_INC_READ;
		ELSIF (SRAM_DATA = '1' AND IO_WRITE = '1') THEN
			STATE <= SRAM_WRITE;
		ELSIF (SRAM_INC_DATA = '1' AND IO_WRITE = '1') THEN
			STATE <= SRAM_INC_WRITE;
		ELSIF (SRAM_ADDR_JPOS = '1' AND IO_WRITE = '1') THEN
			STATE <= JUMP_POS;
		ELSIF (SRAM_ADDR_JNEG = '1' AND IO_WRITE = '1') THEN
			STATE <= JUMP_NEG;
		ELSE 
			STATE <= IDLE;
		END IF;
  
		CASE STATE IS
			WHEN READ_LOWER =>
				IO_DATA(15 DOWNTO 0) <= SRAM_ADDR_ALTERA_SYNTHESIZED(15 DOWNTO 0);
			
			WHEN WRITE_LOWER =>
				SRAM_ADDR_ALTERA_SYNTHESIZED(15 DOWNTO 0) <= IO_DATA(15 DOWNTO 0);
			
			WHEN READ_UPPER =>
				IO_DATA(1 DOWNTO 0) <= SRAM_ADDR_ALTERA_SYNTHESIZED(17 DOWNTO 16);
			
			WHEN WRITE_UPPER =>
				SRAM_ADDR_ALTERA_SYNTHESIZED(17 DOWNTO 16) <= IO_DATA(1 DOWNTO 0);
			
			WHEN SRAM_READ =>
				SRAM_OE_N <= '0';
			
			WHEN SRAM_INC_READ =>
				SRAM_OE_N <= '0';
				
			WHEN SRAM_WRITE =>
				SRAM_WE_N <= '0';
				
			WHEN SRAM_INC_WRITE =>
				SRAM_WE_N <= '0';
				
			WHEN OTHERS =>
				SRAM_OE_N <= '1';
				SRAM_WE_N <= '1';
				IO_DATA <= "ZZZZZZZZZZZZZZZZ";
		END CASE;
		
		IF (PREV_STATE = IDLE AND STATE = JUMP_POS) THEN
			SRAM_ADDR_ALTERA_SYNTHESIZED <= STD_LOGIC_VECTOR(UNSIGNED(SRAM_ADDR_ALTERA_SYNTHESIZED) + UNSIGNED(IO_DATA));
		ELSIF (PREV_STATE = IDLE AND STATE = JUMP_NEG) THEN
			SRAM_ADDR_ALTERA_SYNTHESIZED <= STD_LOGIC_VECTOR(UNSIGNED(SRAM_ADDR_ALTERA_SYNTHESIZED) - UNSIGNED(IO_DATA));
		END IF;
		
		IF (PREV_STATE = SRAM_INC_WRITE OR PREV_STATE = SRAM_INC_READ) AND (PREV_STATE /= STATE) THEN
			SRAM_ADDR_ALTERA_SYNTHESIZED <= STD_LOGIC_VECTOR(UNSIGNED(SRAM_ADDR_ALTERA_SYNTHESIZED) + 1);
		END IF;
    
		PREV_STATE <= STATE;
    END IF;
  END PROCESS;
END bdf_type;